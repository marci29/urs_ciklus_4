-- 10. Definirajte multipleksor s 4 ulaza u VHDL-u korištenjem odabirne logike (entitet i arhitektura) 
