-- 25. Za PicoBlaze procesor napisati sljedeći prekidni potprogram. Na svaki zahtjev za prekid potrebno je očitati stanje vanjske jedinice koja je spojena na IN_PORT. 
-- Na dobivenom podatku ispituje se parnost: ako je paran, potrebno je povećati brojač parnih podataka u ScratchPad memoriji na adresi hex (10),
-- a ukoliko je neparan, povećati brojač neparnih podataka koji se nalazi u ScratchPad memoriji na adresi hex (11).
