-- 20. Potrebno je u VHDL-u projektirati 10-bitni brojač s asinkronim resetom. Brojač ima mogućnost brojanja unaprijed i unatrag što kontrolira pomoću priključka UP_DOWN ( 1 – naprijed, 0 –natrag).
-- Brojač ima na ulazu signal VALUE (4 bita) koji definira vrijednost za koju se povećava ili smanjuje. Brojač na ulazu ima priključke ENABLE ( 1-enable, 0-disable).
-- Prilikom pojave asinkronog reseta svi izlazni signali postavljaju se u 0.
