-- 15. Potrebno je u VHDL‐u projektirati 16‐bitni brojač s asinkronim resetom. 
-- Brojač ima mogućnost brojanja unaprijed i unatrag što se kontrolira pomoću priključka UP_DOWN (‘1’ – unaprijed, ‘0’‐ unatrag). 
-- Brojač ima na ulazu signal VALUE širine 4 bita koji definira vrijednost s kojom se brojač uvećava ili smanjuje. 
-- Brojač na ulazu ima priključak ENABLE koji ako je postavljen u '1' omogućuje brojanje dok u drugom slučaju ga zaustavlja. 
-- Prilikom pojave asinkronog reseta svi izlazni signali sklopa se postavljaju u vrijednost '0'.
