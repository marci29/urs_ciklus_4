/* 5. Definiraj mulitpleksor s 4 ulaza (širina ulaza neka je generičke veličine) korištenjem uvjetne logike u VHDL-u. Potrebno je napisati entitet i arhitekturu. */
