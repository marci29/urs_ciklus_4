/* 7. U VHDL-u opisat sklop za izračun pomičnog prosjeka (Moving Average Filter)... Zadnji zadatak na završnom ispitu 2022. */
