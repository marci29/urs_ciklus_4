-- isti kao 6. https://github.com/marci29/urs_ciklus_4/blob/main/zadatak_6.vhd

-- 6. U VHDL-u definirajte 16-bitno brojilo s asinkronim resetom (prilikom reseta brojilo se postavlja u nulu). Potrebno je napisati entitet i arhitekturu.
