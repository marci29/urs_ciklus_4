-- 6. U VHDL-u definirajte 16-bitno brojilo s asinkronim resetom (prilikom reseta brojilo se postavlja u nulu). Potrebno je napisati entitet i arhitekturu.
