-- 26. Napišite dio VHDL koda (potrebno je napisati samo proces) koji služi za spajanje izlaznih vanjskih jedinica na PicoBlaze? Objasnite kako radi?
-- Napisati primjer korištenja vanjske jedinice u assembleru. 
-- Nacrtati shematski spajanje na KCPSM3 procesor.


